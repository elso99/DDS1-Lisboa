-----------------------------------------------------------------------------
-- Vhdl model created by memgen, (c) 2022 Paulo Flores.
-- Version: 1
-- Command: memgen.pl -s 0
-- Seed: -s 0
-----------------------------------------------------------------------------
library ieee;
library UNISIM;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use UNISIM.Vcomponents.all;

-- Set 0   m[0] = -75 + 22 i		 b[0] = 4 + -7 i
-- i:      Xr +    Xi   =>         Yr  +    Yi 	     Yr     +     Yi
-- 0: x=   26 +   16 i  =>   y=  -2298 +   -635 i  (0xFFFFF706 + 0xFFFFFD85 i)
-- 1: x=   41 +   34 i  =>   y=  -6117 +  -2290 i  (0xFFFFE81B + 0xFFFFF70E i)
-- 2: x=  -38 +  -40 i  =>   y=  -2383 +   -133 i  (0xFFFFF6B1 + 0xFFFFFF7B i)
-- 3: x=  -90 +   41 i  =>   y=   3469 +  -5195 i  (0x00000D8D + 0xFFFFEBB5 i)
-- 4: x=   52 +   75 i  =>   y=  -2077 +  -9683 i  (0xFFFFF7E3 + 0xFFFFDA2D i)
-- 5: x=   22 +   21 i  =>   y=  -4185 + -10781 i  (0xFFFFEFA7 + 0xFFFFD5E3 i)
-- 6: x=  -77 +   93 i  =>   y=   -452 + -19457 i  (0xFFFFFE3C + 0xFFFFB3FF i)
-- 7: x=  -37 +  110 i  =>   y=    -93 + -28528 i  (0xFFFFFFA3 + 0xFFFF9090 i)
-- Sol[0]:		           -11 +  -3566 i  (0xFFFFFFF5 + 0xFFFFF212 i)

-- Set 1   m[1] = -27 + 91 i		 b[1] = -46 + -86 i
-- i:      Xr +    Xi   =>         Yr  +    Yi 	     Yr     +     Yi
-- 0: x=  218 + -170 i  =>   y=   9538 +  24342 i  (0x00002542 + 0x00005F16 i)
-- 1: x=  272 +   -7 i  =>   y=   2785 +  49197 i  (0x00000AE1 + 0x0000C02D i)
-- 2: x=  -76 +   60 i  =>   y=   -669 +  40575 i  (0xFFFFFD63 + 0x00009E7F i)
-- 3: x=  334 + -236 i  =>   y=  11743 +  77255 i  (0x00002DDF + 0x00012DC7 i)
-- 4: x=  -62 +  123 i  =>   y=   2178 +  68206 i  (0x00000882 + 0x00010A6E i)
-- 5: x=  315 + -475 i  =>   y=  36852 + 109610 i  (0x00008FF4 + 0x0001AC2A i)
-- 6: x=  467 +  158 i  =>   y=   9819 + 147755 i  (0x0000265B + 0x0002412B i)
-- 7: x=  338 +   95 i  =>   y=  -7998 + 175862 i  (0xFFFFE0C2 + 0x0002AEF6 i)
-- Sol[1]:		          -999 +  21982 i  (0xFFFFFC19 + 0x000055DE i)

-- Set 2   m[2] = 24 + -7 i		 b[2] = 54 + 22 i
-- i:      Xr +    Xi   =>         Yr  +    Yi 	     Yr     +     Yi
-- 0: x=  228 +  318 i  =>   y=   7752 +   6058 i  (0x00001E48 + 0x000017AA i)
-- 1: x=  330 +   -5 i  =>   y=  15691 +   3650 i  (0x00003D4B + 0x00000E42 i)
-- 2: x= -227 +   64 i  =>   y=  10745 +   6797 i  (0x000029F9 + 0x00001A8D i)
-- 3: x=  141 +  332 i  =>   y=  16507 +  13800 i  (0x0000407B + 0x000035E8 i)
-- 4: x=  403 +  -38 i  =>   y=  25967 +  10089 i  (0x0000656F + 0x00002769 i)
-- 5: x= -378 +  139 i  =>   y=  17922 +  16093 i  (0x00004602 + 0x00003EDD i)
-- 6: x=  481 + -273 i  =>   y=  27609 +   6196 i  (0x00006BD9 + 0x00001834 i)
-- 7: x= -357 + -146 i  =>   y=  18073 +   5213 i  (0x00004699 + 0x0000145D i)
-- Sol[2]:		          2259 +    651 i  (0x000008D3 + 0x0000028B i)

-- Set 3   m[3] = -512 + -512 i		 b[3] = 511 + 511 i
-- i:      Xr +    Xi   =>         Yr  +    Yi 	     Yr     +     Yi
-- 0: x= -512 + -512 i  =>   y=    511 + 524799 i  (0x000001FF + 0x000801FF i)
-- 1: x=  511 +  511 i  =>   y=   1022 +   2046 i  (0x000003FE + 0x000007FE i)
-- 2: x=  511 + -512 i  =>   y= -522243 +   3069 i  (0xFFF807FD + 0x00000BFD i)
-- 3: x= -512 +  511 i  =>   y=   2044 +   4092 i  (0x000007FC + 0x00000FFC i)
-- 4: x= -512 + -512 i  =>   y=   2555 + 528891 i  (0x000009FB + 0x000811FB i)
-- 5: x=  511 + -512 i  =>   y= -520710 + 529914 i  (0xFFF80DFA + 0x000815FA i)
-- 6: x= -512 +  511 i  =>   y=   3577 + 530937 i  (0x00000DF9 + 0x000819F9 i)
-- 7: x=  511 +  511 i  =>   y=   4088 +   8184 i  (0x00000FF8 + 0x00001FF8 i)
-- Sol[3]:		           511 +   1023 i  (0x000001FF + 0x000003FF i)



entity MemIN is
  port (
    clk          : in  std_logic;
    addr_memIN   : in  std_logic_vector(8 downto 0);
    Xr, Xi       : out std_logic_vector(15 downto 0)
    );
end MemIN;


architecture GEN0 of MemIN is
   signal ImRe: std_logic_vector(31 downto 0);
begin

  MEM0_DataIN : RAMB16_S36
    generic map (                       -- memory initialization
      INIT_00 => X"FFB3005D001600150034004BFFA60029FFDAFFD800290022001A0010B51604F9",
      INIT_01 => X"00000000000000000000000000000000000000000000000000000000FFDB006E",
      INIT_02 => X"01D3009E013BFE25FFC2007B014EFF14FFB4003C0110FFF900DAFF56E55BD2AA",
      INIT_03 => X"000000000000000000000000000000000000000000000000000000000152005F",
      INIT_04 => X"01E1FEEFFE86008B0193FFDA008D014CFF1D0040014AFFFB00E4013E18F93616",
      INIT_05 => X"00000000000000000000000000000000000000000000000000000000FE9BFF6E",
      INIT_06 => X"FE0001FF01FFFE00FE00FE00FE0001FF01FFFE0001FF01FFFE00FE000000FFFF",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000001FF01FF",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map (
      CLK   => clk,                     -- Clock
      ADDR  => addr_memIN,              -- 10-bit Address Input
      DI    => x"00000000",             -- 32-bit Data Input
      DIP   => x"0",                    -- 4-bit parity Input
      EN    => '1',                     -- RAM Enable Input
      SSR   => '0',                     -- Synchronous Set/Reset Input
      WE    => '0',                     -- Write Enable Input
      DO    => ImRe,                    -- 32-bit Data Output
      DOP   => open                     -- 1-bit parity Output
      );

   Xr <= ImRe(31 downto 16);
   Xi <= ImRe(15 downto 0);

end GEN0;
